
.SUBCKT INPUT_RES VINP VINN OTA1_INP OTA1_INN GND
xr13 OTA1_INP VINP GND  rppolywo_m lr=10e-6 wr=600e-9 multi=1 m=1 series=5 segspace=250e-9
xr14 VINN OTA1_INN GND  rppolywo_m lr=10e-6 wr=600e-9 multi=1 m=1 series=5 segspace=250e-9
.ENDS



.SUBCKT INVD4BWP_LVT i zn vdd vss

x0 zn i vss vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 

x1 zn i vss vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 

x2 zn i vss vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 

x3 zn i vss vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 

x4 zn i vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

x5 zn i vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

x6 zn i vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

x7 zn i vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 
.ENDS

.SUBCKT DFCND4BWP_LVT_stupid d cp q qn vdd vss

x0 net175 net149 vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

x1 q net149 vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

x2 qn net175 vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

x3 qn net175 vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

xmi43 net12 net145 vdd vdd g45p1lvt l=80e-9 w=240e-9 multi=1 nf=1 

x4 net95 net11 vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

xmi6 net9 d net1 vdd g45p1lvt l=80e-9 w=680e-9 multi=1 nf=1 

x5 qn net175 vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

x6 qn net175 vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

x7 net11 cp vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

x8 q net149 vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

x9 net149 cdn vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

xmi44 net12 cdn vdd vdd g45p1lvt l=80e-9 w=240e-9 multi=1 nf=1 

xmi17 net175 net95 net24 vdd g45p1lvt l=80e-9 w=240e-9 multi=1 nf=1 

x10 net149 net24 vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

x11 net145 net9 vdd vdd g45p1lvt l=80e-9 w=360e-9 multi=1 nf=1 

x12 q net149 vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

xmi16 net145 net11 net24 vdd g45p1lvt l=80e-9 w=360e-9 multi=1 nf=1 

x13 net149 net24 vdd vdd g45p1lvt l=80e-9 w=560e-9 multi=1 nf=1 

x14 net149 cdn vdd vdd g45p1lvt l=80e-9 w=560e-9 multi=1 nf=1 

xmi45 net9 net11 net12 vdd g45p1lvt l=80e-9 w=240e-9 multi=1 nf=1 

x15 q net149 vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

xmi7 net1 net95 vdd vdd g45p1lvt l=80e-9 w=680e-9 multi=1 nf=1 

x16 qn net175 vss vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 

x17 q net149 vss vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 

x18 qn net175 vss vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 

x19 net169 cdn vss vss g45n1lvt l=80e-9 w=400e-9 multi=1 nf=1 

xmi4 net128 net11 vss vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 

x20 qn net175 vss vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 

xmi18 net175 net11 net24 vss g45n1lvt l=80e-9 w=240e-9 multi=1 nf=1 

x21 net145 net9 vss vss g45n1lvt l=80e-9 w=300e-9 multi=1 nf=1 

x22 net149 net24 net169 vss g45n1lvt l=80e-9 w=400e-9 multi=1 nf=1 

xmi15 net145 net95 net24 vss g45n1lvt l=80e-9 w=300e-9 multi=1 nf=1 

x23 net175 net149 vss vss g45n1lvt l=80e-9 w=380e-9 multi=1 nf=1 

x24 q net149 vss vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 

x25 net95 net11 vss vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 

x26 net149 net24 net132 vss g45n1lvt l=80e-9 w=400e-9 multi=1 nf=1 

xmi5 net9 d net128 vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 

x27 net11 cp vss vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 

xmi49 net112 cdn vss vss g45n1lvt l=80e-9 w=240e-9 multi=1 nf=1 

x28 net132 cdn vss vss g45n1lvt l=80e-9 w=400e-9 multi=1 nf=1 

xmi48 net96 net145 net112 vss g45n1lvt l=80e-9 w=240e-9 multi=1 nf=1 

x29 q net149 vss vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 

x30 qn net175 vss vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 

x31 q net149 vss vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 

xmi47 net9 net95 net96 vss g45n1lvt l=80e-9 w=240e-9 multi=1 nf=1 
.ENDS

.SUBCKT OTA_XT_MAGICAL gnd ncas vcm vdd vim vip vom vop

xm29 vs vcmon gnd gnd nch_hvt_mac l=120e-9 w=40.5e-6 multi=1 nf=15 

xm5 pcas vcm bias2 gnd g45n1lvt l=120e-9 w=4.8e-6 multi=1 nf=5 

xm30 tail1 nbias_tail gnd gnd g45n1lvt l=120e-9 w=20e-6 multi=1 nf=25 

xm53 vcmop net0108 vs2 gnd g45n1lvt l=120e-9 w=7.2e-6 multi=1 nf=8 

xm12 vcmon vcm vs2 gnd g45n1lvt l=120e-9 w=7.2e-6 multi=1 nf=8 

xm50 vo1p ncas casn gnd g45n1lvt l=120e-9 w=9e-6 multi=1 nf=10 

xm49 vo1m ncas casp gnd g45n1lvt l=120e-9 w=9e-6 multi=1 nf=10 

xm51 ncas ncas nbias_tail gnd g45n1lvt l=120e-9 w=4e-6 multi=1 nf=5 

xm47 nbias_tail vcm bias1 gnd g45n1lvt l=120e-9 w=4.8e-6 multi=1 nf=5 

xm38 bias1 nbias_tail gnd gnd g45n1lvt l=120e-9 w=4e-6 multi=1 nf=5 

xm7 vop vim vs gnd g45n1lvt l=120e-9 w=36e-6 multi=1 nf=15 

xm43 casn vim tail1 gnd g45n1lvt l=120e-9 w=13.5e-6 multi=1 nf=5 

xm10 vom vip vs gnd g45n1lvt l=120e-9 w=36e-6 multi=1 nf=15 

xm40 casp vip tail1 gnd g45n1lvt l=120e-9 w=13.5e-6 multi=1 nf=5 

xm41 vs2 nbias_tail gnd gnd g45n1lvt l=120e-9 w=14.4e-6 multi=1 nf=10 

xm31 bias2 nbias_tail gnd gnd g45n1lvt l=120e-9 w=4e-6 multi=1 nf=5 

xc0 vo1p net096 cfmom_2t nr=26 lr=1.9e-6 w=70e-9 s=70e-9 stm=2 spm=5 multi=1 ftip=140e-9

xc1 vo1m net096 cfmom_2t nr=26 lr=1.9e-6 w=70e-9 s=70e-9 stm=2 spm=5 multi=1 ftip=140e-9

xc4 vcmon vop cfmom_2t nr=36 lr=4.17e-6 w=70e-9 s=70e-9 stm=2 spm=5 multi=1 ftip=140e-9

xc7 net0108 vop cfmom_2t nr=18 lr=1.91e-6 w=70e-9 s=70e-9 stm=2 spm=4 multi=1 ftip=140e-9

xc3 vcmon vom cfmom_2t nr=36 lr=4.17e-6 w=70e-9 s=70e-9 stm=2 spm=5 multi=1 ftip=140e-9

xc6 net0108 vom cfmom_2t nr=18 lr=1.91e-6 w=70e-9 s=70e-9 stm=2 spm=4 multi=1 ftip=140e-9
xr10 net0108 vom gnd  rppolywo_m lr=3.6e-6 wr=400e-9 multi=1 m=1 series=6 segspace=250e-9

xr1 vop net0108 gnd  rppolywo_m lr=3.6e-6 wr=400e-9 multi=1 m=1 series=6 segspace=250e-9

xr8 vo1m net096 gnd  rppolywo_m lr=7.86e-6 wr=400e-9 multi=1 m=1 series=10 segspace=250e-9

xr2 net096 vo1p gnd  rppolywo_m lr=7.86e-6 wr=400e-9 multi=1 m=1 series=10 segspace=250e-9


xm57 vo1p pcas cas2n vdd g45p1lvt l=120e-9 w=18e-6 multi=1 nf=10 

xm64 vcmon vcmop vdd vdd g45p1lvt l=120e-9 w=9.6e-6 multi=1 nf=10 

xm67 vom vo1p vdd vdd g45p1lvt l=120e-9 w=28.8e-6 multi=1 nf=20 

xm66 vcmop vcmop vdd vdd g45p1lvt l=120e-9 w=9.6e-6 multi=1 nf=10 

xm8 cas2n net096 vdd vdd g45p1lvt l=120e-9 w=12e-6 multi=1 nf=10 

xm61 cas2p net096 vdd vdd g45p1lvt l=120e-9 w=12e-6 multi=1 nf=10 

xm56 vo1m pcas cas2p vdd g45p1lvt l=120e-9 w=18e-6 multi=1 nf=10 

xm9 vop vo1m vdd vdd g45p1lvt l=120e-9 w=28.8e-6 multi=1 nf=20 

xm58 pcas pcas net088 vdd g45p1lvt l=120e-9 w=6.4e-6 multi=1 nf=4 

xm63 net088 pcas vdd vdd pch_hvt_mac l=120e-9 w=1.07e-6 multi=1 nf=1 
.ENDS

.SUBCKT OTA_XT_MAGICAL_2 gnd ncas vcm vdd vim vip vom vop

xm29 vs vcmon gnd gnd nch_hvt_mac l=120e-9 w=40.5e-6 multi=1 nf=20 

xm5 pcas vcm bias2 gnd g45n1lvt l=120e-9 w=4.8e-6 multi=1 nf=5 

xm30 tail1 nbias_tail gnd gnd g45n1lvt l=120e-9 w=20e-6 multi=1 nf=25 

xm53 vcmop net0108 vs2 gnd g45n1lvt l=120e-9 w=7.2e-6 multi=1 nf=8 

xm12 vcmon vcm vs2 gnd g45n1lvt l=120e-9 w=7.2e-6 multi=1 nf=8 

xm50 vo1p ncas casn gnd g45n1lvt l=120e-9 w=9e-6 multi=1 nf=10 

xm49 vo1m ncas casp gnd g45n1lvt l=120e-9 w=9e-6 multi=1 nf=10 

xm51 ncas ncas nbias_tail gnd g45n1lvt l=120e-9 w=4e-6 multi=1 nf=5 

xm47 nbias_tail vcm bias1 gnd g45n1lvt l=120e-9 w=4.8e-6 multi=1 nf=5 

xm38 bias1 nbias_tail gnd gnd g45n1lvt l=120e-9 w=4e-6 multi=1 nf=5 

xm7 vop vim vs gnd g45n1lvt l=120e-9 w=36e-6 multi=1 nf=15 

xm43 casn vim tail1 gnd g45n1lvt l=120e-9 w=13.5e-6 multi=1 nf=5 

xm10 vom vip vs gnd g45n1lvt l=120e-9 w=36e-6 multi=1 nf=15 

xm40 casp vip tail1 gnd g45n1lvt l=120e-9 w=13.5e-6 multi=1 nf=5 

xm41 vs2 nbias_tail gnd gnd g45n1lvt l=120e-9 w=14.4e-6 multi=1 nf=10 

xm31 bias2 nbias_tail gnd gnd g45n1lvt l=120e-9 w=4e-6 multi=1 nf=5 

xc0 vo1p net096 cfmom_2t nr=26 lr=1.9e-6 w=70e-9 s=70e-9 stm=2 spm=5 multi=1 ftip=140e-9

xc1 vo1m net096 cfmom_2t nr=26 lr=1.9e-6 w=70e-9 s=70e-9 stm=2 spm=5 multi=1 ftip=140e-9

xc4 vcmon vop cfmom_2t nr=36 lr=4.17e-6 w=70e-9 s=70e-9 stm=2 spm=5 multi=1 ftip=140e-9

xc7 net0108 vop cfmom_2t nr=18 lr=1.91e-6 w=70e-9 s=70e-9 stm=2 spm=4 multi=1 ftip=140e-9

xc3 vcmon vom cfmom_2t nr=36 lr=4.17e-6 w=70e-9 s=70e-9 stm=2 spm=5 multi=1 ftip=140e-9

xc6 net0108 vom cfmom_2t nr=18 lr=1.91e-6 w=70e-9 s=70e-9 stm=2 spm=4 multi=1 ftip=140e-9
xr10 net0108 vom gnd  rppolywo_m lr=3.6e-6 wr=400e-9 multi=1 m=1 series=6 segspace=250e-9

xr1 vop net0108 gnd  rppolywo_m lr=3.6e-6 wr=400e-9 multi=1 m=1 series=6 segspace=250e-9

xr8 vo1m net096 gnd  rppolywo_m lr=7.86e-6 wr=400e-9 multi=1 m=1 series=10 segspace=250e-9

xr2 net096 vo1p gnd  rppolywo_m lr=7.86e-6 wr=400e-9 multi=1 m=1 series=10 segspace=250e-9


xm57 vo1p pcas cas2n vdd g45p1lvt l=120e-9 w=18e-6 multi=1 nf=10 

xm64 vcmon vcmop vdd vdd g45p1lvt l=120e-9 w=9.6e-6 multi=1 nf=10 

xm67 vom vo1p vdd vdd g45p1lvt l=120e-9 w=28.8e-6 multi=1 nf=20 

xm66 vcmop vcmop vdd vdd g45p1lvt l=120e-9 w=9.6e-6 multi=1 nf=10 

xm8 cas2n net096 vdd vdd g45p1lvt l=120e-9 w=12e-6 multi=1 nf=10 

xm61 cas2p net096 vdd vdd g45p1lvt l=120e-9 w=12e-6 multi=1 nf=10 

xm56 vo1m pcas cas2p vdd g45p1lvt l=120e-9 w=18e-6 multi=1 nf=10 

xm9 vop vo1m vdd vdd g45p1lvt l=120e-9 w=28.8e-6 multi=1 nf=20 

xm58 pcas pcas net088 vdd g45p1lvt l=120e-9 w=6.4e-6 multi=1 nf=4 

xm63 net088 pcas vdd vdd pch_hvt_mac l=120e-9 w=1.07e-6 multi=1 nf=1 
.ENDS



.SUBCKT BUFFD4BWP_LVT i z vdd vss

x0 z net11 vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

x1 net11 i vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

x2 net11 i vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

x3 z net11 vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

x4 z net11 vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

x5 z net11 vdd vdd g45p1lvt l=80e-9 w=820e-9 multi=1 nf=1 

x6 z net11 vss vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 

x7 z net11 vss vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 

x8 z net11 vss vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 

x9 net11 i vss vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 

x10 z net11 vss vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 

x11 net11 i vss vss g45n1lvt l=80e-9 w=620e-9 multi=1 nf=1 
.ENDS

.SUBCKT NR2D8BWP_LVT a1 a2 zn vdd vss

x0 net13 a2 vdd vdd g45p1lvt l=80e-9 w=6.56e-6 multi=1 nf=1 

x1 zn a1 net13 vdd g45p1lvt l=80e-9 w=6.56e-6 multi=1 nf=1 

x2 zn a2 vss vss g45n1lvt l=80e-9 w=4.96e-6 multi=1 nf=1 

x3 zn a1 vss vss g45n1lvt l=80e-9 w=4.96e-6 multi=1 nf=1 
.ENDS

.SUBCKT SR_Latch_LVT q qb r s vdd vss


xi1 r qb q vdd vss NR2D8BWP_LVT


xi0 s q qb vdd vss NR2D8BWP_LVT
.ENDS

.SUBCKT COMPARATOR_schematic clk gnd outm outp vdd _net0 _net1

xm0 gnd intern gnd gnd g45n1lvt l=1e-6 w=1.05e-6 multi=1 nf=1 

xm22 gnd interp gnd gnd g45n1lvt l=1e-6 w=1.05e-6 multi=1 nf=1 

xm16 outm crossp gnd gnd g45n1lvt l=40e-9 w=1.44e-6 multi=1 nf=4 

xm17 outp crossn gnd gnd g45n1lvt l=40e-9 w=1.44e-6 multi=1 nf=4 

xm4 crossn crossp intern gnd g45n1lvt l=40e-9 w=1.92e-6 multi=1 nf=4 

xm3 crossp crossn interp gnd g45n1lvt l=40e-9 w=1.92e-6 multi=1 nf=4 

xm7 net069 clk gnd gnd g45n1lvt l=40e-9 w=3.68e-6 multi=1 nf=8 

xm5 intern _net0 net069 gnd g45n1lvt l=40e-9 w=7.68e-6 multi=1 nf=8 

xm6 interp _net1 net069 gnd g45n1lvt l=40e-9 w=7.68e-6 multi=1 nf=8 

xm8 outm crossp vdd vdd g45p1lvt l=40e-9 w=1.92e-6 multi=1 nf=4 

xm18 intern clk vdd vdd g45p1lvt l=40e-9 w=960e-9 multi=1 nf=2 

xm15 outp crossn vdd vdd g45p1lvt l=40e-9 w=1.92e-6 multi=1 nf=4 

xm2 interp clk vdd vdd g45p1lvt l=40e-9 w=960e-9 multi=1 nf=2 

xm1 crossn clk vdd vdd g45p1lvt l=40e-9 w=960e-9 multi=1 nf=2 

xm12 crossp clk vdd vdd g45p1lvt l=40e-9 w=960e-9 multi=1 nf=2 

xm14 crossn crossp vdd vdd g45p1lvt l=40e-9 w=3.84e-6 multi=1 nf=8 

xm13 crossp crossn vdd vdd g45p1lvt l=40e-9 w=3.84e-6 multi=1 nf=8 
.ENDS

.SUBCKT RR1 net040 net010 VREF GND net025 SYS_CLKB VDD net035
xi24 net040 net010 VREF GND BUFFD4BWP_LVT
xi25 net025 SYS_CLKB net040 net035 VDD GND DFCND4BWP_LVT_stupid
.ENDS

.SUBCKT RRR1 net046 SYS_CLKB VDD DO net038 GND net025 net028 net020 SYS_CLK
xi12 net046 SYS_CLKB DO net038 VDD GND DFCND4BWP_LVT_stupid
xi6 net046 net025 net028 net020 VDD GND SR_Latch_LVT
xi4 SYS_CLK SYS_CLKB VDD GND INVD4BWP_LVT
.ENDS

.SUBCKT GPDK_CDL_TEST DO GND IBIAS1 IBIAS2 SYS_CLK VCM VDD VINN VINP OTA1_INN OTA1_INP OTA2_INN OTA2_INP SUM_N SUM_P VINT1N VINT1P VINT2N VINT2P VREF

input_res  VINP VINN OTA1_INP OTA1_INN GND INPUT_RES

xr47 OTA1_INN VINT2P GND  rppolywo_m lr=34.8e-6 wr=400e-9 multi=1 m=1 series=46 segspace=250e-9

xr28 OTA1_INP VINT2N GND  rppolywo_m lr=34.8e-6 wr=400e-9 multi=1 m=1 series=46 segspace=250e-9

xr21 net010 OTA1_INP GND  rppolywo_m lr=10e-6 wr=600e-9 multi=1 m=1 series=5 segspace=250e-9

xr20 net012 OTA1_INN GND  rppolywo_m lr=10e-6 wr=600e-9 multi=1 m=1 series=5 segspace=250e-9

xr23 net010 OTA2_INP GND  rppolywo_m lr=10e-6 wr=600e-9 multi=1 m=1 series=10 segspace=250e-9

xr25 net012 SUM_N GND  rppolywo_m lr=10e-6 wr=600e-9 multi=1 m=1 series=15 segspace=250e-9

xr24 net010 SUM_P GND  rppolywo_m lr=10e-6 wr=600e-9 multi=1 m=1 series=15 segspace=250e-9

xr22 net012 OTA2_INN GND  rppolywo_m lr=10e-6 wr=600e-9 multi=1 m=1 series=10 segspace=250e-9

xr19 VINT2N SUM_N GND   rppolywo_m lr=10e-6 wr=600e-9 multi=1 m=1 series=1 segspace=250e-9

xr16 VINT1N OTA2_INN GND  rppolywo_m lr=10e-6 wr=600e-9 multi=1 m=1 series=5 segspace=250e-9

xr17 VINT1P OTA2_INP GND  rppolywo_m lr=10e-6 wr=600e-9 multi=1 m=1 series=5 segspace=250e-9


xr18  VINT2P SUM_P GND   rppolywo_m lr=10e-6 wr=600e-9 multi=1 m=1 series=1 segspace=250e-9




xc4 OTA1_INP VINT1N cfmom_2t nr=96 lr=12.4e-6 w=70e-9 s=70e-9 stm=2 spm=5 multi=1 ftip=140e-9

xc2 OTA2_INN VINT2P cfmom_2t nr=70 lr=9.85e-6 w=70e-9 s=70e-9 stm=2 spm=5 multi=1 ftip=140e-9

xc0 OTA1_INN VINT1P cfmom_2t nr=96 lr=12.4e-6 w=70e-9 s=70e-9 stm=2 spm=5 multi=1 ftip=140e-9

xc1 OTA2_INP VINT2N cfmom_2t nr=70 lr=9.85e-6 w=70e-9 s=70e-9 stm=2 spm=5 multi=1 ftip=140e-9








xi22 GND IBIAS2 VCM VDD OTA2_INN OTA2_INP VINT2N VINT2P OTA_XT_MAGICAL


xi20 GND IBIAS1 VCM VDD OTA1_INP OTA1_INN VINT1P VINT1N OTA_XT_MAGICAL








xi19 SYS_CLK GND net028 net020 VDD SUM_P SUM_N COMPARATOR_schematic

rr1 net040 net010 VREF GND net025 SYS_CLKB VDD net035 RR1
rr2 net026 net012 VREF GND net046 SYS_CLKB VDD net022 RR1


rrr1 net046 SYS_CLKB VDD DO net038 GND net025 net028 net020 SYS_CLK RRR1

.ENDS
